// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Thu Oct 05 14:13:55 2023
//
// Verilog Description of module main
//

module main (CK, DAC1A, DAC1B, DAC1C, DAC1D, DAC1E, DAC1F, DAC1G, 
            DAC1H, DAC2A, DAC2B, DAC2C, DAC2D, DAC2E, DAC2F, DAC2G, 
            DAC2H, A, B, C, D, E, F, G, H, K, L, M, 
            N, O, P, Q, R, S, T, V, W, UPLOAD, EMPTY, 
            ACTIV);   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(10[8:12])
    input CK;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(12[3:5])
    output DAC1A;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(14[3:8])
    output DAC1B;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(15[3:8])
    output DAC1C;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(16[3:8])
    output DAC1D;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(17[3:8])
    output DAC1E;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(18[3:8])
    output DAC1F;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(19[3:8])
    output DAC1G;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(20[3:8])
    output DAC1H;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(21[3:8])
    output DAC2A;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(22[3:8])
    output DAC2B;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(23[3:8])
    output DAC2C;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(24[3:8])
    output DAC2D;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(25[3:8])
    output DAC2E;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(26[3:8])
    output DAC2F;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(27[3:8])
    output DAC2G;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(28[3:8])
    output DAC2H;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(29[3:8])
    output A;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(30[3:4])
    output B;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(31[3:4])
    output C;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(32[3:4])
    output D;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(33[3:4])
    output E;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(34[3:4])
    output F;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(35[3:4])
    output G;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(36[3:4])
    output H;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(37[3:4])
    output K;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(38[3:4])
    output L;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(39[3:4])
    output M;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(40[3:4])
    output N;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(41[3:4])
    output O;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(42[3:4])
    output P;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(43[3:4])
    output Q;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(44[3:4])
    output R;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(45[3:4])
    output S;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(46[3:4])
    output T;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(47[3:4])
    output V;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(48[3:4])
    output W;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(49[3:4])
    output UPLOAD;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(50[3:9])
    output EMPTY;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(51[3:8])
    output ACTIV;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(52[3:8])
    
    wire CK_c /* synthesis is_clock=1, SET_AS_NETWORK=CK_c */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(12[3:5])
    
    wire GND_net, VCC_net, n138, L_c, n137;
    wire [12:0]\Clock_Divider.count ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(91[11:16])
    wire [12:0]\Clock_Divider.count_12__N_14 ;
    
    wire n140, n136, n135, n134;
    wire [12:0]\Clock_Divider.count_12__N_1 ;
    
    wire n133, L_N_28, n24, n13, n21, n20, n17, n20_adj_1, n17_adj_2, 
        n16, n177;
    
    VHI i2 (.Z(VCC_net));
    OB M_pad (.I(VCC_net), .O(M));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(40[3:4])
    FD1S3AX SCK_15 (.D(L_N_28), .CK(CK_c), .Q(L_c));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam SCK_15.GSR = "ENABLED";
    CCU2D add_7_9 (.A0(\Clock_Divider.count [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n136), .COUT(n137), .S0(\Clock_Divider.count_12__N_14 [7]), 
          .S1(\Clock_Divider.count_12__N_14 [8]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(\Clock_Divider.count [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n137), .COUT(n138), .S0(\Clock_Divider.count_12__N_14 [9]), 
          .S1(\Clock_Divider.count_12__N_14 [10]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    FD1S3AX \Clock_Divider.count_i1  (.D(\Clock_Divider.count_12__N_1 [1]), 
            .CK(CK_c), .Q(\Clock_Divider.count [1]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i1 .GSR = "ENABLED";
    OB L_pad (.I(L_c), .O(L));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(39[3:4])
    OB DAC1B_pad (.I(GND_net), .O(DAC1B));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(15[3:8])
    OB K_pad (.I(GND_net), .O(K));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(38[3:4])
    LUT4 i94_4_lut_rep_1 (.A(\Clock_Divider.count [7]), .B(n24), .C(n20), 
         .D(\Clock_Divider.count [6]), .Z(n177)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i94_4_lut_rep_1.init = 16'h0001;
    OB H_pad (.I(VCC_net), .O(H));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(37[3:4])
    OB G_pad (.I(VCC_net), .O(G));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(36[3:4])
    OB F_pad (.I(GND_net), .O(F));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(35[3:4])
    OB E_pad (.I(VCC_net), .O(E));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(34[3:4])
    OB D_pad (.I(VCC_net), .O(D));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(33[3:4])
    OB C_pad (.I(GND_net), .O(C));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(32[3:4])
    OB B_pad (.I(VCC_net), .O(B));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(31[3:4])
    OB A_pad (.I(VCC_net), .O(A));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(30[3:4])
    OB DAC2H_pad (.I(GND_net), .O(DAC2H));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(29[3:8])
    OB DAC2G_pad (.I(GND_net), .O(DAC2G));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(28[3:8])
    OB DAC2F_pad (.I(GND_net), .O(DAC2F));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(27[3:8])
    OB DAC2E_pad (.I(GND_net), .O(DAC2E));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(26[3:8])
    OB DAC2D_pad (.I(GND_net), .O(DAC2D));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(25[3:8])
    OB DAC2C_pad (.I(GND_net), .O(DAC2C));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(24[3:8])
    OB DAC2B_pad (.I(GND_net), .O(DAC2B));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(23[3:8])
    OB DAC2A_pad (.I(GND_net), .O(DAC2A));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(22[3:8])
    OB DAC1H_pad (.I(GND_net), .O(DAC1H));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(21[3:8])
    OB DAC1G_pad (.I(GND_net), .O(DAC1G));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(20[3:8])
    OB DAC1F_pad (.I(GND_net), .O(DAC1F));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(19[3:8])
    OB DAC1E_pad (.I(GND_net), .O(DAC1E));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(18[3:8])
    OB DAC1D_pad (.I(GND_net), .O(DAC1D));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(17[3:8])
    OB DAC1C_pad (.I(GND_net), .O(DAC1C));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(16[3:8])
    LUT4 i2_2_lut (.A(\Clock_Divider.count_12__N_14 [5]), .B(\Clock_Divider.count_12__N_14 [6]), 
         .Z(n13)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(121[6:26])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i9_4_lut (.A(n17_adj_2), .B(n13), .C(\Clock_Divider.count_12__N_14 [11]), 
         .D(\Clock_Divider.count_12__N_14 [2]), .Z(n20_adj_1)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(121[6:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i72_2_lut_2_lut (.A(n177), .B(\Clock_Divider.count_12__N_14 [1]), 
         .Z(\Clock_Divider.count_12__N_1 [1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i72_2_lut_2_lut.init = 16'h4444;
    VLO i1 (.Z(GND_net));
    OB DAC1A_pad (.I(CK_c), .O(DAC1A));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(14[3:8])
    OB N_pad (.I(VCC_net), .O(N));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(41[3:4])
    OB O_pad (.I(GND_net), .O(O));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(42[3:4])
    OB P_pad (.I(VCC_net), .O(P));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(43[3:4])
    OB Q_pad (.I(VCC_net), .O(Q));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(44[3:4])
    OB R_pad (.I(VCC_net), .O(R));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(45[3:4])
    OB S_pad (.I(GND_net), .O(S));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(46[3:4])
    OB T_pad (.I(VCC_net), .O(T));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(47[3:4])
    OB V_pad (.I(GND_net), .O(V));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(48[3:4])
    OB W_pad (.I(CK_c), .O(W));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(49[3:4])
    OB UPLOAD_pad (.I(GND_net), .O(UPLOAD));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(50[3:9])
    OB EMPTY_pad (.I(GND_net), .O(EMPTY));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(51[3:8])
    OB ACTIV_pad (.I(GND_net), .O(ACTIV));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(52[3:8])
    IB CK_pad (.I(CK), .O(CK_c));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(12[3:5])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i4_2_lut (.A(\Clock_Divider.count [1]), .B(\Clock_Divider.count [0]), 
         .Z(n17)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i71_2_lut_2_lut (.A(n177), .B(\Clock_Divider.count_12__N_14 [0]), 
         .Z(\Clock_Divider.count_12__N_1 [0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i71_2_lut_2_lut.init = 16'h4444;
    CCU2D add_7_13 (.A0(\Clock_Divider.count [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n138), .S0(\Clock_Divider.count_12__N_14 [11]), 
          .S1(\Clock_Divider.count_12__N_14 [12]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(\Clock_Divider.count [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n135), .COUT(n136), .S0(\Clock_Divider.count_12__N_14 [5]), 
          .S1(\Clock_Divider.count_12__N_14 [6]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(\Clock_Divider.count [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n134), .COUT(n135), .S0(\Clock_Divider.count_12__N_14 [3]), 
          .S1(\Clock_Divider.count_12__N_14 [4]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(\Clock_Divider.count [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\Clock_Divider.count [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n133), .COUT(n134), .S0(\Clock_Divider.count_12__N_14 [1]), 
          .S1(\Clock_Divider.count_12__N_14 [2]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\Clock_Divider.count [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n133), .S1(\Clock_Divider.count_12__N_14 [0]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(117[14:19])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    TSALL TSALL_INST (.TSALL(GND_net));
    FD1S3IX \Clock_Divider.count_i3  (.D(\Clock_Divider.count_12__N_14 [3]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [3]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i3 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i4  (.D(\Clock_Divider.count_12__N_14 [4]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [4]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i4 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i5  (.D(\Clock_Divider.count_12__N_14 [5]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [5]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i5 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i6  (.D(\Clock_Divider.count_12__N_14 [6]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [6]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i6 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i7  (.D(\Clock_Divider.count_12__N_14 [7]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [7]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i7 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i8  (.D(\Clock_Divider.count_12__N_14 [8]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [8]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i8 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i9  (.D(\Clock_Divider.count_12__N_14 [9]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [9]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i9 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i10  (.D(\Clock_Divider.count_12__N_14 [10]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [10]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i10 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i11  (.D(\Clock_Divider.count_12__N_14 [11]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [11]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i11 .GSR = "ENABLED";
    FD1S3IX \Clock_Divider.count_i12  (.D(\Clock_Divider.count_12__N_14 [12]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [12]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i12 .GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut (.A(n177), .B(\Clock_Divider.count_12__N_14 [1]), 
         .C(n140), .D(\Clock_Divider.count_12__N_14 [0]), .Z(L_N_28)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i1_4_lut_4_lut.init = 16'h5450;
    LUT4 i6_3_lut (.A(\Clock_Divider.count_12__N_14 [8]), .B(\Clock_Divider.count_12__N_14 [7]), 
         .C(\Clock_Divider.count_12__N_14 [3]), .Z(n17_adj_2)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(121[6:26])
    defparam i6_3_lut.init = 16'hfefe;
    FD1S3IX \Clock_Divider.count_i2  (.D(\Clock_Divider.count_12__N_14 [2]), 
            .CK(CK_c), .CD(n177), .Q(\Clock_Divider.count [2]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i2 .GSR = "ENABLED";
    LUT4 i7_3_lut (.A(\Clock_Divider.count [10]), .B(\Clock_Divider.count [8]), 
         .C(\Clock_Divider.count [3]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i5_2_lut (.A(\Clock_Divider.count_12__N_14 [10]), .B(\Clock_Divider.count_12__N_14 [12]), 
         .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(121[6:26])
    defparam i5_2_lut.init = 16'heeee;
    FD1S3AX \Clock_Divider.count_i0  (.D(\Clock_Divider.count_12__N_1 [0]), 
            .CK(CK_c), .Q(\Clock_Divider.count [0]));   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(98[2] 126[9])
    defparam \Clock_Divider.count_i0 .GSR = "ENABLED";
    LUT4 i8_4_lut (.A(\Clock_Divider.count [12]), .B(\Clock_Divider.count [4]), 
         .C(\Clock_Divider.count [5]), .D(\Clock_Divider.count [9]), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i8_4_lut.init = 16'hfffe;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i11_4_lut (.A(n21), .B(n17), .C(\Clock_Divider.count [11]), .D(\Clock_Divider.count [2]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(114[7:26])
    defparam i11_4_lut.init = 16'hfeff;
    LUT4 i10_4_lut (.A(\Clock_Divider.count_12__N_14 [4]), .B(n20_adj_1), 
         .C(n16), .D(\Clock_Divider.count_12__N_14 [9]), .Z(n140)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/nathan sayer/documents/osi/kicad/a305001a (function generator)/p3050fg/main.vhd(121[6:26])
    defparam i10_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

